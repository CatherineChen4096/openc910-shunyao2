module TOP();

	top ();
endmodule 
