module TOP();

	top_top ();
endmodule 

module top_top();
    top ();
endmodule
